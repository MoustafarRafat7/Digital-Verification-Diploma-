interface shift_reg_interface ();

bit reset, serial_in, direction, mode; 
bit [5:0] datain, dataout;


endinterface