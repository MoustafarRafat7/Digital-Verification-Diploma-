package Memory_Package;

parameter T = 2;

class Memory_Transaction;

rand logic [7:0] DATA_IN;
rand logic [15:0] ADDRESS;

endclass

endpackage